module log_x_map (
    input  logic        clk,
    input  logic        rst,
    
    input  logic [9:0]  pixel_x,    // 0-799
    input  logic        active,
    
    output logic [8:0]  bin_index,  // 0-511
    output logic        bin_valid
);

    
    logic [8:0] lut [0:799] = '{
    9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0,
    9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0,
    9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0,
    9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0,
    9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0,
    9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0,
    9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0,
    9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0,
    9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0,
    9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0,
    9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0, 9'd  0,
    9'd  0, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1,
    9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1,
    9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1,
    9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1,
    9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1,
    9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1,
    9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  1, 9'd  2, 9'd  2, 9'd  2,
    9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2,
    9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2,
    9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2,
    9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2, 9'd  2,
    9'd  2, 9'd  2, 9'd  3, 9'd  3, 9'd  3, 9'd  3, 9'd  3, 9'd  3,
    9'd  3, 9'd  3, 9'd  3, 9'd  3, 9'd  3, 9'd  3, 9'd  3, 9'd  3,
    9'd  3, 9'd  3, 9'd  3, 9'd  3, 9'd  3, 9'd  3, 9'd  3, 9'd  3,
    9'd  3, 9'd  3, 9'd  3, 9'd  3, 9'd  3, 9'd  3, 9'd  3, 9'd  4,
    9'd  4, 9'd  4, 9'd  4, 9'd  4, 9'd  4, 9'd  4, 9'd  4, 9'd  4,
    9'd  4, 9'd  4, 9'd  4, 9'd  4, 9'd  4, 9'd  4, 9'd  4, 9'd  4,
    9'd  4, 9'd  4, 9'd  4, 9'd  4, 9'd  4, 9'd  4, 9'd  5, 9'd  5,
    9'd  5, 9'd  5, 9'd  5, 9'd  5, 9'd  5, 9'd  5, 9'd  5, 9'd  5,
    9'd  5, 9'd  5, 9'd  5, 9'd  5, 9'd  5, 9'd  5, 9'd  5, 9'd  5,
    9'd  5, 9'd  5, 9'd  6, 9'd  6, 9'd  6, 9'd  6, 9'd  6, 9'd  6,
    9'd  6, 9'd  6, 9'd  6, 9'd  6, 9'd  6, 9'd  6, 9'd  6, 9'd  6,
    9'd  6, 9'd  6, 9'd  6, 9'd  7, 9'd  7, 9'd  7, 9'd  7, 9'd  7,
    9'd  7, 9'd  7, 9'd  7, 9'd  7, 9'd  7, 9'd  7, 9'd  7, 9'd  7,
    9'd  7, 9'd  7, 9'd  8, 9'd  8, 9'd  8, 9'd  8, 9'd  8, 9'd  8,
    9'd  8, 9'd  8, 9'd  8, 9'd  8, 9'd  8, 9'd  8, 9'd  8, 9'd  9,
    9'd  9, 9'd  9, 9'd  9, 9'd  9, 9'd  9, 9'd  9, 9'd  9, 9'd  9,
    9'd  9, 9'd  9, 9'd  9, 9'd  9, 9'd 10, 9'd 10, 9'd 10, 9'd 10,
    9'd 10, 9'd 10, 9'd 10, 9'd 10, 9'd 10, 9'd 10, 9'd 10, 9'd 11,
    9'd 11, 9'd 11, 9'd 11, 9'd 11, 9'd 11, 9'd 11, 9'd 11, 9'd 11,
    9'd 11, 9'd 12, 9'd 12, 9'd 12, 9'd 12, 9'd 12, 9'd 12, 9'd 12,
    9'd 12, 9'd 12, 9'd 12, 9'd 13, 9'd 13, 9'd 13, 9'd 13, 9'd 13,
    9'd 13, 9'd 13, 9'd 13, 9'd 14, 9'd 14, 9'd 14, 9'd 14, 9'd 14,
    9'd 14, 9'd 14, 9'd 14, 9'd 14, 9'd 15, 9'd 15, 9'd 15, 9'd 15,
    9'd 15, 9'd 15, 9'd 15, 9'd 16, 9'd 16, 9'd 16, 9'd 16, 9'd 16,
    9'd 16, 9'd 16, 9'd 16, 9'd 17, 9'd 17, 9'd 17, 9'd 17, 9'd 17,
    9'd 17, 9'd 17, 9'd 18, 9'd 18, 9'd 18, 9'd 18, 9'd 18, 9'd 18,
    9'd 19, 9'd 19, 9'd 19, 9'd 19, 9'd 19, 9'd 19, 9'd 20, 9'd 20,
    9'd 20, 9'd 20, 9'd 20, 9'd 20, 9'd 21, 9'd 21, 9'd 21, 9'd 21,
    9'd 21, 9'd 21, 9'd 22, 9'd 22, 9'd 22, 9'd 22, 9'd 22, 9'd 22,
    9'd 23, 9'd 23, 9'd 23, 9'd 23, 9'd 23, 9'd 24, 9'd 24, 9'd 24,
    9'd 24, 9'd 24, 9'd 25, 9'd 25, 9'd 25, 9'd 25, 9'd 25, 9'd 26,
    9'd 26, 9'd 26, 9'd 26, 9'd 27, 9'd 27, 9'd 27, 9'd 27, 9'd 27,
    9'd 28, 9'd 28, 9'd 28, 9'd 28, 9'd 29, 9'd 29, 9'd 29, 9'd 29,
    9'd 30, 9'd 30, 9'd 30, 9'd 30, 9'd 31, 9'd 31, 9'd 31, 9'd 31,
    9'd 32, 9'd 32, 9'd 32, 9'd 32, 9'd 33, 9'd 33, 9'd 33, 9'd 33,
    9'd 34, 9'd 34, 9'd 34, 9'd 35, 9'd 35, 9'd 35, 9'd 35, 9'd 36,
    9'd 36, 9'd 36, 9'd 37, 9'd 37, 9'd 37, 9'd 37, 9'd 38, 9'd 38,
    9'd 38, 9'd 39, 9'd 39, 9'd 39, 9'd 40, 9'd 40, 9'd 40, 9'd 41,
    9'd 41, 9'd 41, 9'd 42, 9'd 42, 9'd 42, 9'd 43, 9'd 43, 9'd 43,
    9'd 44, 9'd 44, 9'd 44, 9'd 45, 9'd 45, 9'd 45, 9'd 46, 9'd 46,
    9'd 47, 9'd 47, 9'd 47, 9'd 48, 9'd 48, 9'd 48, 9'd 49, 9'd 49,
    9'd 50, 9'd 50, 9'd 50, 9'd 51, 9'd 51, 9'd 52, 9'd 52, 9'd 53,
    9'd 53, 9'd 53, 9'd 54, 9'd 54, 9'd 55, 9'd 55, 9'd 56, 9'd 56,
    9'd 56, 9'd 57, 9'd 57, 9'd 58, 9'd 58, 9'd 59, 9'd 59, 9'd 60,
    9'd 60, 9'd 61, 9'd 61, 9'd 62, 9'd 62, 9'd 63, 9'd 63, 9'd 64,
    9'd 64, 9'd 65, 9'd 65, 9'd 66, 9'd 66, 9'd 67, 9'd 67, 9'd 68,
    9'd 68, 9'd 69, 9'd 70, 9'd 70, 9'd 71, 9'd 71, 9'd 72, 9'd 72,
    9'd 73, 9'd 74, 9'd 74, 9'd 75, 9'd 75, 9'd 76, 9'd 76, 9'd 77,
    9'd 78, 9'd 78, 9'd 79, 9'd 80, 9'd 80, 9'd 81, 9'd 82, 9'd 82,
    9'd 83, 9'd 83, 9'd 84, 9'd 85, 9'd 86, 9'd 86, 9'd 87, 9'd 88,
    9'd 88, 9'd 89, 9'd 90, 9'd 90, 9'd 91, 9'd 92, 9'd 93, 9'd 93,
    9'd 94, 9'd 95, 9'd 96, 9'd 96, 9'd 97, 9'd 98, 9'd 99, 9'd 99,
    9'd100, 9'd101, 9'd102, 9'd103, 9'd103, 9'd104, 9'd105, 9'd106,
    9'd107, 9'd108, 9'd108, 9'd109, 9'd110, 9'd111, 9'd112, 9'd113,
    9'd114, 9'd115, 9'd116, 9'd116, 9'd117, 9'd118, 9'd119, 9'd120,
    9'd121, 9'd122, 9'd123, 9'd124, 9'd125, 9'd126, 9'd127, 9'd128,
    9'd129, 9'd130, 9'd131, 9'd132, 9'd133, 9'd134, 9'd135, 9'd136,
    9'd137, 9'd139, 9'd140, 9'd141, 9'd142, 9'd143, 9'd144, 9'd145,
    9'd146, 9'd148, 9'd149, 9'd150, 9'd151, 9'd152, 9'd154, 9'd155,
    9'd156, 9'd157, 9'd158, 9'd160, 9'd161, 9'd162, 9'd164, 9'd165,
    9'd166, 9'd167, 9'd169, 9'd170, 9'd171, 9'd173, 9'd174, 9'd176,
    9'd177, 9'd178, 9'd180, 9'd181, 9'd183, 9'd184, 9'd186, 9'd187,
    9'd188, 9'd190, 9'd191, 9'd193, 9'd194, 9'd196, 9'd198, 9'd199,
    9'd201, 9'd202, 9'd204, 9'd205, 9'd207, 9'd209, 9'd210, 9'd212,
    9'd214, 9'd215, 9'd217, 9'd219, 9'd221, 9'd222, 9'd224, 9'd226,
    9'd228, 9'd229, 9'd231, 9'd233, 9'd235, 9'd237, 9'd239, 9'd240,
    9'd242, 9'd244, 9'd246, 9'd248, 9'd250, 9'd252, 9'd254, 9'd256,
    9'd258, 9'd260, 9'd262, 9'd264, 9'd266, 9'd268, 9'd271, 9'd273,
    9'd275, 9'd277, 9'd279, 9'd281, 9'd284, 9'd286, 9'd288, 9'd290,
    9'd293, 9'd295, 9'd297, 9'd300, 9'd302, 9'd304, 9'd307, 9'd309,
    9'd312, 9'd314, 9'd317, 9'd319, 9'd322, 9'd324, 9'd327, 9'd329,
    9'd332, 9'd334, 9'd337, 9'd340, 9'd342, 9'd345, 9'd348, 9'd350,
    9'd353, 9'd356, 9'd359, 9'd362, 9'd364, 9'd367, 9'd370, 9'd373,
    9'd376, 9'd379, 9'd382, 9'd385, 9'd388, 9'd391, 9'd394, 9'd397,
    9'd400, 9'd404, 9'd407, 9'd410, 9'd413, 9'd416, 9'd420, 9'd423,
    9'd426, 9'd430, 9'd433, 9'd436, 9'd440, 9'd443, 9'd447, 9'd450,
    9'd454, 9'd457, 9'd461, 9'd465, 9'd468, 9'd472, 9'd476, 9'd479,
    9'd483, 9'd487, 9'd491, 9'd495, 9'd499, 9'd503, 9'd507, 9'd511
};

    always_ff @(posedge clk) begin
        if (rst) begin
            bin_index <= '0;
            bin_valid <= 1'b0;
        end else begin
            bin_index <= lut[pixel_x];
            bin_valid <= active;
        end
    end

endmodule